module kitten

// square calculates the second power of `x`
pub fn square(x int) int {
	return x * x
}
